`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.02.2020 13:05:30
// Design Name: 
// Module Name: test_clk_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_clk_tb(
    );
  reg           clk_50m;  
  reg   [10:0]  sw;
  reg   [4:0]   btn;
  wire  [9:0]   led;
  wire  [6:0]   hex0;
  wire  [6:0]   hex1;
  wire  [6:0]   hex2;
  wire  [6:0]   hex3;
  wire  [7:0]   hex_on;
    
  mainframe DUT (
  .clk_50m (  clk_50m  ),
  .sw      (  sw       ),
  .btn     (  btn      ),
  .led     (  led      ),
  .hex0    (  hex0     ),
  .hex1    (  hex1     ),
  .hex2    (  hex2     ),
  .hex3    (  hex3     ),
  .hex_on  (  hex_on   )
  );

 initial begin
    //��������� ���� � ����������� ������� debounce
    sw[10:0] = 11'b00000000000;
    btn[4:0] = 5'b11111;
    #50;
    
    //��������� ����� �� key_3
    btn[4]=1'b0;
    #100;
    btn[4]=1'b1;
    
    #200;
    
    //���������� ������������� (���� ��)
    sw[10:0] = 11'b00000000111;
    
    #200
    
    //������ ������ � ������� �� key_0
    btn[0]=1'b0;
    #100;
    btn[0]=1'b1;
    
    #200;
    
    btn[1]=1'b0;
    #100;
    btn[1]=1'b1;
    
    #200
    
    //������ ������ � ������� �� key_0 (��� ��������� ��������� ������
    btn[0]=1'b0;
    #100;
    btn[0]=1'b1;
    
    #200;
    
    btn[1]=1'b0;
    #100;
    btn[1]=1'b1;
    
    #200
    
    sw[10:0] = 11'b00000000011;
    
    #200;
    
    btn[0]=1'b0;
    #100;
    btn[0]=1'b1;
    
    #200;
    
    btn[1]=1'b0;
    #100;
    btn[1]=1'b1;
    
    #200
    
    btn[4]=1'b0;
    #100;
    btn[4]=1'b1;   
 
    //��������� ���� � ���������� ������� debounce
//    sw[10:0] = 11'b10000000000;
//    btn[4:0] = 5'b11111;
//    #50;
    
//    //��������� ����� �� key_3
//    btn[4]=1'b0;
//    #100;
//    btn[4]=1'b1;
    
//    #200;
    
//    //���������� ������������� (���� ��)
//    sw[10:0] = 11'b10000000111;
    
//    #200
    
//    //������ ������ � ������� �� key_0
//    btn[0]=1'b0;
//    #150;
//    btn[0]=1'b1;
    
//    #200;
    
//    //������ ������ � ������� �� key_0 (��� ��������� ��������� ������
//    btn[0]=1'b0;
//    #150;
//    btn[0]=1'b1;
    
//    #200;
    
//    sw[10:0] = 11'b10000000011;
    
//    #200;
    
//    btn[0]=1'b0;
//    #150;
//    btn[0]=1'b1;
    
//    #200;
    
//    btn[4]=1'b0;
//    #150;
//    btn[4]=1'b1;   
 end 
 
 //��������� CLK �������
 always begin //�������� 1-0 CLK �������
    clk_50m = 1'b1;
    #10;
    clk_50m = 1'b0;
    #10;
 end
    
endmodule
