module counter(
    input [9:0] SW,
    input [1:0] KEY,
    output [9:0] LEDR,
    output [6:0] HEX1,
    output [6:0] HEX0
);

 /*
    You shall add your code here
  */

endmodule