module counter(
    input clk100_i,
    input rstn_i,
    input [9:0] sw_i,
    input [1:0] key_i,
    output [9:0] ledr_o,
    output [6:0] hex1_o,
    output [6:0] hex0_o
);

// Haaaaaaands

endmodule