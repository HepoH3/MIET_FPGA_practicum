`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.05.2020 18:33:32
// Design Name: 
// Module Name: mainframe
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//������ mainframe
//�� ��� ����������, ������ ��� ��� �� �������.
//������� - ��� Counter_10
module mainframe(                           
  input      [10:0]  sw_i,                    //���� ��������������
  //��������!!! sw[10] ������������ ��� ��������� ������� "debounce" ��� ������. �������� ������ = 1 
  input      [4:0]  btn_i,                    //���� ������ (btn[0]=key0, btn[4]=key1, btn[1]=key2)
  input             clk_50m,                //���� ��������� ������� �������� 50 ���
  output     [9:0]  ledr_o,                    //����� �� ���������� 
  output     [6:0]  hex0_o,                   //����� �� ������ �������������� ���������
  output     [6:0]  hex1_o,                   //����� �� ������ �������������� ���������
  output     [6:0]  hex2_o,                   //����� �� ������ �������������� ���������
  output     [6:0]  hex3_o,                   //����� �� �������� �������������� ���������
  output     [7:0]  hex_on_o                  //����� ������������� ��������������� ���������� �� 8 (0 - ��������)
    );
     
  wire  [9:0]  register;              //���� �������� (��������� �������� ���������� ��������������)
  wire  [7:0]  counter_1;             //���� ������� �������� (������� ������������ �� ����� ����� ���������� ������. � �������)
  wire  [7:0]  counter_2;             //���� ������� �������� (������� ������������ �� ����� ����� ���������� ������. � �������)
  assign ledr_o   = register;          //���������� �������� � ������ �� ����������
  assign hex_on_o = 8'b1111_0000;      //�������� ������ 4 ���������������
  
  //����/����� �������� �� ������ hub
  hub u1(                         
    .btn_i        (  btn_i[4:0]      ),
    .sw_i         (  sw_i[10:0]      ),
    .clk_50m      (  clk_50m         ),
    .register_o   (  register[9:0]   ),
    .counter_1_o  (  counter_1[7:0]  ),
    .counter_2_o  (  counter_2[7:0]  )
  );
  
  //����������� ������ �� �������������� ����������:
  //������ �������
  decoder_8 u2 (
    .bit4_0_i     (  counter_1[3:0]  ),
    .bit4_1_i     (  counter_1[7:4]  ),
    .segment_0_o  (  hex0_o[6:0]     ),
    .segment_1_o  (  hex1_o[6:0]     )
  );
  //������ �������
  decoder_8 u3 (
    .bit4_0_i     (  counter_2[3:0]  ),
    .bit4_1_i     (  counter_2[7:4]  ),
    .segment_0_o  (  hex2_o[6:0]     ),
    .segment_1_o  (  hex3_o[6:0]     )
  );
endmodule
