`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.05.2020 18:33:32
// Design Name: 
// Module Name: mainframe
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//������ mainframe (������� - "mainfr")
module mainframe(                           
  input      [9:0]  sw,                     //���� ��������������
  input      [4:0]  btn,                    //���� ������ 
  input             clk_50m,               //���� ��������� ������� �������� 50 ���
  output     [9:0]  led,                    //����� �� ���������� 
  output reg [6:0]  hex,                    //����� �� ��������� �������������� ���������
  output reg [7:0]  hex_on                  //����� ������������� ��������������� ���������� �� 8 (0 - ��������)
    );
     
  wire [9:0]register;                //���� �������� (��������� �������� ���������� ��������������)
  wire [7:0]counter;                 //���� �������� (������� ������������ �� ����� ����� ���������� ������. � �������)
  assign led = register;             //���������� �������� � ������ �� ����������
  
  //����/����� �������� �� ������ KEY_Switching (������� - "KS")
  hub u1(                         
    .btn_i(btn[4:0]),
    .sw_i(sw[9:0]),
    .clk_50m(clk_50m),
    .register_o(register[9:0]),
    .counter_o(counter[7:0])
  );
  
  //���������� ������ �� �������������� ����������:
  //��� ������ ����������� ��������, ���������������� 0-1-0... � �������� clk_50m, ���������� ������������ ����� ����� ������������
  reg disp_selector = 1'd0;          //���������� ������� ������
  always @(posedge clk_50m) begin          //�������� ���������� �� 0->1 
      disp_selector <= disp_selector + 1'b1; 
      if (disp_selector == 1'b0)
      begin
          hex_on <= 8'b1111_1110;
          case (counter[3:0])        //�� ������ ��������� ��������� ������ 4 ���� ��������
              4'd0  : hex = 7'b100_0000;
              4'd1  : hex = 7'b111_1001;
              4'd2  : hex = 7'b010_0100;
              4'd3  : hex = 7'b011_0000;
              4'd4  : hex = 7'b001_1001;
              4'd5  : hex = 7'b001_0010;
              4'd6  : hex = 7'b000_0010;
              4'd7  : hex = 7'b111_1000;
              4'd8  : hex = 7'b000_0000;
              4'd9  : hex = 7'b001_0000;
              4'd10 : hex = 7'b000_1000;
              4'd11 : hex = 7'b000_0011;
              4'd12 : hex = 7'b100_0110;
              4'd13 : hex = 7'b010_0001;
              4'd14 : hex = 7'b000_0110;
              4'd15 : hex = 7'b000_1110;
          endcase
      end
      
      if (disp_selector == 1'b1)
      begin
          hex_on <= 8'b1111_1101;
          case (counter[7:4])        //�� ������ ��������� ��������� ������ 4 ���� ��������
              4'd0  : hex = 7'b100_0000;
              4'd1  : hex = 7'b111_1001;
              4'd2  : hex = 7'b010_0100;
              4'd3  : hex = 7'b011_0000;
              4'd4  : hex = 7'b001_1001;
              4'd5  : hex = 7'b001_0010;
              4'd6  : hex = 7'b000_0010;
              4'd7  : hex = 7'b111_1000;
              4'd8  : hex = 7'b000_0000;
              4'd9  : hex = 7'b001_0000;
              4'd10 : hex = 7'b000_1000;
              4'd11 : hex = 7'b000_0011;
              4'd12 : hex = 7'b100_0110;
              4'd13 : hex = 7'b010_0001;
              4'd14 : hex = 7'b000_0110;
              4'd15 : hex = 7'b000_1110;
          endcase
      end    
  end
  
endmodule
